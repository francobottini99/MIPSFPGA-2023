`ifndef __IS_ZERO_VH__
`define __IS_ZERO_VH__
    `include "common.vh"

    `define DEFAULT_IS_ZERO_BUS_SIZE `ARQUITECTURE_BITS
`endif // __IS_ZERO_VH__