`ifndef __MEM_VH__
`define __MEM_VH__
    `include "data_memory.vh"

    `define DEFAULT_MEM_BUS_SIZE `ARQUITECTURE_BITS 
`endif // __MEM_VH__