`ifndef __IS_NOT_EQUAL_VH__
`define __IS_NOT_EQUAL_VH__
    `include "common.vh"

    `define DEFAULT_IS_NOT_EQUAL_BUS_SIZE `ARQUITECTURE_BITS
`endif // __IS_NOT_EQUAL_VH__