`ifndef __ID_EX_VH__
`define __ID_EX_VH__
    `include "id.vh"
    `include "ex.vh"
`endif // __ID_EX_VH__