`ifndef __ALU_CONTROL_VH__
`define __ALU_CONTROL_VH__
    `include "common.vh"
    `include "codes.vh"

    `define DEFAULT_ALU_OP_BUS_WIDTH    6
    `define DEFAULT_ALU_FUNCT_BUS_WIDTH 6
    `define DEFAULT_ALU_CTR_BUS_WIDTH   4
`endif // __ALU_CONTROL_VH__