`ifndef __ALU_VH__
`define __ALU_VH__
    `include "common.vh"
    `include "alu_control.vh"
    
    `define DEFAULT_ALU_IO_BUS_WIDTH  8
`endif // __ALU_VH__