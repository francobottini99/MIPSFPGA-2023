`ifndef __UART_VH__
`define __UART_VH__
    `define DEFAULT_UART_DATA_BITS 8
    `define DEFAULT_UART_SB_TICKS  16
    `define DEFAULT_UART_DVSR_BIT  9
    `define DEFAULT_UART_DVSR      326
    `define DEFAULT_UART_FIFO_SIZE 8
`endif // __UART_VH__