`ifndef __SHIFT_LEFT_VH__
`define __SHIFT_LEFT_VH__
    `include "common.vh"

    `define DEFAULT_SHIFT_LEFT_BUS_SIZE `ARQUITECTURE_BITS
    `define DEFAULT_SHIFT_LEFT          2
`endif // __SHIFT_LEFT_VH__