`ifndef __WB_VH__
`define __WB_VH__
    `include "common.vh"

    `define DEFAULT_WB_IO_BUS_SIZE `ARQUITECTURE_BITS 
`endif // __WB_VH__