`ifndef __SHORT_CIRCUIT_VH__
`define __SHORT_CIRCUIT_VH__
    `include "common.vh"
    `include "codes.vh"

    `define DEFAULT_SHORT_CIRCUIT_MEM_ADDR_SIZE 5
`endif // __SHORT_CIRCUIT_VH__