`timescale 1ns / 1ps

`include "tb.vh"
`include "codes.vh"

module tb_main_control;

    reg           i_bus_a_not_equal_bus_b;
    reg           i_instruction_is_nop;
    reg  [5 : 0]  i_op;
    reg  [5 : 0]  i_funct;
    wire [19 : 0] o_ctrl_regs;

    main_control dut 
    (
        .i_bus_a_not_equal_bus_b (i_bus_a_not_equal_bus_b),
        .i_instruction_is_nop    (i_instruction_is_nop),
        .i_op                    (i_op),
        .i_funct                 (i_funct),
        .o_ctrl_regs             (o_ctrl_regs)
    );

    initial 
    begin
        i_instruction_is_nop = `LOW;
        
        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_ADD;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST ADD  ERROR");
        else
            $display("TEST ADD  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SUB;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SUB  ERROR");
        else
            $display("TEST SUB  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_AND;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST AND  ERROR");
        else
            $display("TEST AND  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_OR;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST OR   ERROR");
        else
            $display("TEST OR   PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_XOR;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST XOR  ERROR");
        else
            $display("TEST XOR  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_NOR;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST NOR  ERROR");
        else
            $display("TEST NOR  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SLT;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SLT  ERROR");
        else
            $display("TEST SLT  PASS");
        
        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SLL;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_SHAMT, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SLL  ERROR");
        else
            $display("TEST SLL  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SRL;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_SHAMT, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SRL  ERROR");
        else
            $display("TEST SRL  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SRA;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_SHAMT, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SRA  ERROR");
        else
            $display("TEST SRA  PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_ADDU;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST ADDU ERROR");
        else
            $display("TEST ADDU PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SUBU;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SUBU ERROR");
        else
            $display("TEST SUBU PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SLLV;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SLLV ERROR");
        else
            $display("TEST SLLV PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SRLV;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SRLV ERROR");
        else
            $display("TEST SRLV PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_SRAV;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RD, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_BUS_B, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SRAV ERROR");
        else
            $display("TEST SRAV PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_JALR;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_NOT_SEQ, `CODE_MAIN_CTR_JMP_REG, `CODE_MAIN_CTR_REG_DST_GPR_31, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_NEXT_SEQ_PC, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE,  `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST JALR ERROR");
        else
            $display("TEST JALR PASS");

        i_op    = `CODE_OP_R_TYPE;
        i_funct = `CODE_FUNCT_JR;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_NOT_SEQ, `CODE_MAIN_CTR_JMP_REG, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NOTHING, `CODE_ALU_CTR_R_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST JR   ERROR");
        else
            $display("TEST JR   PASS");
            
        i_funct = 0;
        
        i_op = `CODE_OP_LW;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_WORD, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_MEM_RESULT }))
            $display("TEST LW   ERROR");
        else
            $display("TEST LW   PASS");
        
        i_op = `CODE_OP_SW;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_BUS_A, `CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_STORE_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_WORD, `CODE_MAIN_CTR_MEM_WRITE_ENABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST SW   ERROR");
        else
            $display("TEST SW   PASS");

        i_op = `CODE_OP_BEQ;
        i_bus_a_not_equal_bus_b = `HIGH;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NOTHING, `CODE_ALU_CTR_BRANCH_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST BEQ1 ERROR");
        else
            $display("TEST BEQ1 PASS");

        i_op = `CODE_OP_BEQ;
        i_bus_a_not_equal_bus_b = `LOW;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_NOT_SEQ, `CODE_MAIN_CTR_JMP_BRANCH, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NOTHING, `CODE_ALU_CTR_BRANCH_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST BEQ2 ERROR");
        else
            $display("TEST BEQ2 PASS");

        i_op = `CODE_OP_BNE;
        i_bus_a_not_equal_bus_b = `LOW;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NOTHING, `CODE_ALU_CTR_BRANCH_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST BNE1 ERROR");
        else
            $display("TEST BNE1 PASS");

        i_op = `CODE_OP_BNE;
        i_bus_a_not_equal_bus_b = `HIGH;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_NOT_SEQ, `CODE_MAIN_CTR_JMP_BRANCH, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NOTHING, `CODE_ALU_CTR_BRANCH_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST BNE2 ERROR");
        else
            $display("TEST BNE2 PASS");

        i_op = `CODE_OP_ADDI;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_ADDI, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST ADDI ERROR");
        else
            $display("TEST ADDI PASS");

        i_op = `CODE_OP_J;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_NOT_SEQ, `CODE_MAIN_CTR_JMP_DIR, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NOTHING, `CODE_ALU_CTR_JUMP_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST J    ERROR");
        else
            $display("TEST J    PASS");

        i_op = `CODE_OP_JAL;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_NOT_SEQ, `CODE_MAIN_CTR_JMP_DIR, `CODE_MAIN_CTR_REG_DST_GPR_31, `CODE_ALU_CTR_SRC_A_NOTHING, `CODE_ALU_CTR_SRC_B_NEXT_SEQ_PC, `CODE_ALU_CTR_JUMP_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST JAL  ERROR");
        else
            $display("TEST JAL  PASS");

        i_op = `CODE_OP_ANDI;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_USIG_INM,  `CODE_ALU_CTR_ANDI, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST ANDI ERROR");
        else
            $display("TEST ANDI PASS");
        
        i_op = `CODE_OP_ORI;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_USIG_INM,  `CODE_ALU_CTR_ORI, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST ORI  ERROR");
        else
            $display("TEST ORI  PASS");

        i_op = `CODE_OP_XORI;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_USIG_INM,  `CODE_ALU_CTR_XORI, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST XORI ERROR");
        else
            $display("TEST XORI PASS");

        i_op = `CODE_OP_SLTI;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_SLTI, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST SLTI ERROR");
        else
            $display("TEST SLTI PASS");

        i_op = `CODE_OP_LUI;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_UPPER_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_ALU_RESULT }))
            $display("TEST LUI  ERROR");
        else
            $display("TEST LUI  PASS");

        i_op = `CODE_OP_LB;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_SIG_BYTE, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_MEM_RESULT }))
            $display("TEST LB   ERROR");
        else
            $display("TEST LB   PASS");

        i_op = `CODE_OP_LBU;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_USIG_BYTE, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_MEM_RESULT }))
            $display("TEST LBU  ERROR");
        else
            $display("TEST LBU  PASS");

        i_op = `CODE_OP_LH;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_SIG_HALFWORD, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_MEM_RESULT }))
            $display("TEST LH   ERROR");
        else
            $display("TEST LH   PASS");

        i_op = `CODE_OP_LHU;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_USIG_HALFWORD, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_MEM_RESULT }))
            $display("TEST LHU  ERROR");
        else
            $display("TEST LHU  PASS");

        i_op = `CODE_OP_LWU;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_RT, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_LOAD_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_WORD, `CODE_MAIN_CTR_MEM_WR_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WRITE_DISABLE, `CODE_MAIN_CTR_WB_ENABLE, `CODE_MAIN_CTR_MEM_TO_REG_MEM_RESULT }))
            $display("TEST LWU  ERROR");
        else
            $display("TEST LWU  PASS");

        i_op = `CODE_OP_SB;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_STORE_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_BYTE, `CODE_MAIN_CTR_MEM_WRITE_ENABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST SB   ERROR");
        else
            $display("TEST SB   PASS");

        i_op = `CODE_OP_SH;
        #10;
        if (!(o_ctrl_regs === { `CODE_MAIN_CTR_NEXT_PC_SRC_SEQ, `CODE_MAIN_CTR_NOT_JMP, `CODE_MAIN_CTR_REG_DST_NOTHING, `CODE_ALU_CTR_SRC_A_BUS_A,`CODE_ALU_CTR_SRC_B_SIG_INM, `CODE_ALU_CTR_STORE_TYPE, `CODE_MAIN_CTR_MEM_RD_SRC_NOTHING, `CODE_MAIN_CTR_MEM_WR_SRC_HALFWORD, `CODE_MAIN_CTR_MEM_WRITE_ENABLE, `CODE_MAIN_CTR_WB_DISABLE, `CODE_MAIN_CTR_MEM_TO_REG_NOTHING }))
            $display("TEST SH   ERROR");
        else
            $display("TEST SH   PASS");
        
        $finish;
    end

endmodule