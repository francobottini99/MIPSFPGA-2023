`ifndef __DEBUGGER_CONTROL_VH__
`define __DEBUGGER_CONTROL_VH__
    `include "common.vh"

    `define DEFAULT_DEBUGGER_CONTROL_UART_BUS_SIZE           8
    `define DEFAULT_DEBUGGER_CONTROL_OUT_BUS_SIZE           `DEFAULT_DEBUGGER_CONTROL_UART_BUS_SIZE * 7
    `define DEFAULT_DEBUGGER_CONTROL_IN_BUS_SIZE            `DEFAULT_DEBUGGER_CONTROL_UART_BUS_SIZE * 4
    `define DEFAULT_DEBUGGER_CONTROL_REGISTER_SIZE          `ARQUITECTURE_BITS

    `define DEBUGGER_CONTROL_STATE_WAIT_RD                      5'b00000
    `define DEBUGGER_CONTROL_STATE_WAIT_RD_TRANSITION           5'b00001
    `define DEBUGGER_CONTROL_STATE_WAIT_WR                      5'b00010
    `define DEBUGGER_CONTROL_STATE_WAIT_WR_TRANSITION           5'b00011 
    `define DEBUGGER_CONTROL_STATE_UNKNOWN_CMD                  5'b00100
    `define DEBUGGER_CONTROL_STATE_END_PROGRAM                  5'b00101
    `define DEBUGGER_CONTROL_STATE_EMPTY_PROGRAM                5'b00110
    `define DEBUGGER_CONTROL_STATE_END_STEP                     5'b00111
    `define DEBUGGER_CONTROL_STATE_DECODE                       5'b01000
    `define DEBUGGER_CONTROL_STATE_IDLE                         5'b01001
    `define DEBUGGER_CONTROL_STATE_FLUSH                        5'b01010
    `define DEBUGGER_CONTROL_STATE_RESET                        5'b01011
    `define DEBUGGER_CONTROL_STATE_LOAD_IDLE                    5'b01100
    `define DEBUGGER_CONTROL_STATE_LOAD                         5'b01101
    `define DEBUGGER_CONTROL_STATE_RUN_DECODE                   5'b01110
    `define DEBUGGER_CONTROL_STATE_RUN_WAIT_TRANSITION          5'b01111
    `define DEBUGGER_CONTROL_STATE_RUN_IDLE                     5'b10000
    `define DEBUGGER_CONTROL_STATE_RUN_BY_STEPS                 5'b10001
    `define DEBUGGER_CONTROL_STATE_RUN                          5'b10010
    `define DEBUGGER_CONTROL_STATE_PRINT_REGISTERS_TRANSITION   5'b10011
    `define DEBUGGER_CONTROL_STATE_PRINT_REGISTERS              5'b10100
    `define DEBUGGER_CONTROL_STATE_PRINT_MEMORY_DATA_TRANSITION 5'b10101
    `define DEBUGGER_CONTROL_STATE_PRINT_MEMORY_DATA            5'b10110

`endif // __DEBUGGER_CONTROL_VH__