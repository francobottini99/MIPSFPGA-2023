`ifndef __INSTRUCTION_MEMORY_VH__
`define __INSTRUCTION_MEMORY_VH__
    `include "common.vh"

    `define DEFAULT_INSTRUCTION_MEMORY_WORD_SIZE_IN_BYTES `ARQUITECTURE_BITS / `BYTE_SIZE 
    `define DEFAULT_INSTRUCTION_MEMORY_MEM_SIZE_IN_WORDS  10
    `define DEFAULT_INSTRUCTION_MEMORY_PC_SIZE            `ARQUITECTURE_BITS
`endif // __INSTRUCTION_MEMORY_VH__