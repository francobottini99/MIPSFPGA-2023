`ifndef __MEMORY_PRINTER_VH__
`define __MEMORY_PRINTER_VH__
    `include "common.vh"

    `define DEFAULT_MEMORY_PRINTER_UART_BUS_SIZE        8
    `define DEFAULT_MEMORY_PRINTER_OUT_BUS_SIZE         `DEFAULT_MEMORY_PRINTER_UART_BUS_SIZE * 7
    `define DEFAULT_MEMORY_PRINTER_MEMORY_SLOT_SIZE     `ARQUITECTURE_BITS
    `define DEFAULT_MEMORY_PRINTER_MEMORY_DATA_BUS_SIZE `DEFAULT_MEMORY_PRINTER_MEMORY_SLOT_SIZE * 32

    `define MEMORY_PRINTER_STATE_IDLE               2'b00
    `define MEMORY_PRINTER_STATE_PRINT              2'b01
    `define MEMORY_PRINTER_STATE_WAIT_WR_TRANSITION 2'b10
    `define MEMORY_PRINTER_STATE_WAIT_WR            2'b11

`endif // __MEMORY_PRINTER_VH__