`ifndef __EX_MEM_VH__
`define __EX_MEM_VH__
    `include "ex.vh"
    `include "mem.vh"
`endif // __EX_MEM_VH__