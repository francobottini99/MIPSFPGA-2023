`ifndef __IF_VH__
`define __IF_VH__
    `include "pc.vh"
    `include "instruction_memory.vh"
`endif // __IF_VH__