`ifndef __EX_VH__
`define __EX_VH__
    `include "alu.vh"
    `include "alu_control.vh"

    `define DEFAULT_EX_BUS_SIZE `ARQUITECTURE_BITS
`endif // __EX_VH__