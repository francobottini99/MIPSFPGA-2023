`ifndef __SIG_EXTEND_VH__
`define __SIG_EXTEND_VH__
    `include "common.vh"
    
    `define DEFAULT_SIG_EXTEND_OUT_REG_SIZE `ARQUITECTURE_BITS
    `define DEFAULT_SIG_EXTEND_IN_REG_SIZE  16
`endif // __SIG_EXTEND_VH__