`ifndef __MEM_WB_VH__
`define __MEM_WB_VH__
    `include "mem.vh"
    `include "wb.vh"
`endif // __MEM_WB_VH__