`ifndef __UNSIG_EXTEND_VH__
`define __UNSIG_EXTEND_VH__
    `include "common.vh"
    
    `define DEFAULT_UNSIG_EXTEND_OUT_REG_SIZE `ARQUITECTURE_BITS
    `define DEFAULT_UNSIG_EXTEND_IN_REG_SIZE  16
`endif // __UNSIG_EXTEND_VH__