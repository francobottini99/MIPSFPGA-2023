`ifndef __ADDER_VH__
`define __ADDER_VH__
    `include "common.vh"

    `define DEFAULT_ADDER_BUS_SIZE `ARQUITECTURE_BITS
`endif // __ADDER_VH__