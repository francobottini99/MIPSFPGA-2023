`ifndef __RISK_DETECTION_VH__
`define __RISK_DETECTION_VH__
    `include "common.vh"
    `include "codes.vh"
`endif // __RISK_DETECTION_VH__