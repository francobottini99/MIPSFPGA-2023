`ifndef __MAIN_CONTROL_VH__
`define __MAIN_CONTROL_VH__
    `include "common.vh"
    `include "codes.vh"
`endif // __MAIN_CONTROL_VH__