`ifndef __DATA_MEMORY_VH__
`define __DATA_MEMORY_VH__
    `include "common.vh"

    `define DEFAULT_DATA_MEMORY_ADDR_SIZE 5
    `define DEFAULT_DATA_MEMORY_SLOT_SIZE `ARQUITECTURE_BITS
`endif // __DATA_MEMORY_VH__