`ifndef __REGISTERS_BANK_VH__
`define __REGISTERS_BANK_VH__
    `include "common.vh"
    
    `define DEFAULT_REGISTERS_BANK_SIZE 32
    `define DEFAULT_REGISTERS_SIZE      32
`endif // __REGISTERS_BANK_VH__