`ifndef __UART_BRG_VH__
`define __UART_BRG_VH__    
    `define BAUDRATE_PRECISION 4
    `define BAUDRATE_PERIOD    10
`endif // __UART_BRG_VH__