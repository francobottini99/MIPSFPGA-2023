`ifndef __MIPS_VH__
`define __MIPS_VH__
    `include "common.vh"
    `include "if.vh"
    `include "id.vh"
    `include "ex.vh"
    `include "mem.vh"
    `include "wb.vh"
`endif // __MIPS_VH__