`ifndef __IF_ID_VH__
`define __IF_ID_VH__
    `include "if.vh"
    `include "id.vh"
`endif // __IF_ID_VH__