`ifndef __MUX_VH__
`define __MUX_VH__
    `include "common.vh"

    `define DEFAULT_MUX_CHANNELS 2
    `define DEFAULT_MUX_BUS_SIZE `ARQUITECTURE_BITS
`endif // __MUX_VH__